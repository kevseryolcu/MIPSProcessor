library verilog;
use verilog.vl_types.all;
entity or32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end or32Bit;
