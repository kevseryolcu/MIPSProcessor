library verilog;
use verilog.vl_types.all;
entity nor32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end nor32Bit;
