library verilog;
use verilog.vl_types.all;
entity xor32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end xor32Bit;
