library verilog;
use verilog.vl_types.all;
entity fullAdder16Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end fullAdder16Bit;
