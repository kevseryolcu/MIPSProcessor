library verilog;
use verilog.vl_types.all;
entity ALU32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end ALU32Bit;
