library verilog;
use verilog.vl_types.all;
entity mux8to1 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end mux8to1;
