module mux8to1for32Bit(S[2:0], I0[31:0], I1[31:0], I2[31:0], I3[31:0], I4[31:0], I5[31:0], I6[31:0], I7[31:0], Result[31:0]);
	input [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
	input [2:0] S;
	output [31:0] Result;
	
	mux8to1 g0(Result[0], S, I0[0], I1[0], I2[0], I3[0], I4[0], I5[0], I6[0], I7[0]);
	mux8to1 g1(Result[1], S, I0[1], I1[1], I2[1], I3[1], I4[1], I5[1], I6[1], I7[1]);
	mux8to1 g2(Result[2], S, I0[2], I1[2], I2[2], I3[2], I4[2], I5[2], I6[2], I7[2]);
	mux8to1 g3(Result[3], S, I0[3], I1[3], I2[3], I3[3], I4[3], I5[3], I6[3], I7[3]);
	mux8to1 g4(Result[4], S, I0[4], I1[4], I2[4], I3[4], I4[4], I5[4], I6[4], I7[4]);
	mux8to1 g5(Result[5], S, I0[5], I1[5], I2[5], I3[5], I4[5], I5[5], I6[5], I7[5]);
	mux8to1 g6(Result[6], S, I0[6], I1[6], I2[6], I3[6], I4[6], I5[6], I6[6], I7[6]);
	mux8to1 g7(Result[7], S, I0[7], I1[7], I2[7], I3[7], I4[7], I5[7], I6[7], I7[7]);
	mux8to1 g8(Result[8], S, I0[8], I1[8], I2[8], I3[8], I4[8], I5[8], I6[8], I7[8]);
	mux8to1 g9(Result[9], S, I0[9], I1[9], I2[9], I3[9], I4[9], I5[9], I6[9], I7[9]);
	mux8to1 g10(Result[10], S, I0[10], I1[10], I2[10], I3[10], I4[10], I5[10], I6[10], I7[10]);
	mux8to1 g11(Result[11], S, I0[11], I1[11], I2[11], I3[11], I4[11], I5[11], I6[11], I7[11]);
	mux8to1 g12(Result[12], S, I0[12], I1[12], I2[12], I3[12], I4[12], I5[12], I6[12], I7[12]);
	mux8to1 g13(Result[13], S, I0[13], I1[13], I2[13], I3[13], I4[13], I5[13], I6[13], I7[13]);
	mux8to1 g14(Result[14], S, I0[14], I1[14], I2[14], I3[14], I4[14], I5[14], I6[14], I7[14]);
	mux8to1 g15(Result[15], S, I0[15], I1[15], I2[15], I3[15], I4[15], I5[15], I6[15], I7[15]);
	mux8to1 g16(Result[16], S, I0[16], I1[16], I2[16], I3[16], I4[16], I5[16], I6[16], I7[16]);
	mux8to1 g17(Result[17], S, I0[17], I1[17], I2[17], I3[17], I4[17], I5[17], I6[17], I7[17]);
	mux8to1 g18(Result[18], S, I0[18], I1[18], I2[18], I3[18], I4[18], I5[18], I6[18], I7[18]);
	mux8to1 g19(Result[19], S, I0[19], I1[19], I2[19], I3[19], I4[19], I5[19], I6[19], I7[19]);
	mux8to1 g20(Result[20], S, I0[20], I1[20], I2[20], I3[20], I4[20], I5[20], I6[20], I7[20]);
	mux8to1 g21(Result[21], S, I0[21], I1[21], I2[21], I3[21], I4[21], I5[21], I6[21], I7[21]);
	mux8to1 g22(Result[22], S, I0[22], I1[22], I2[22], I3[22], I4[22], I5[22], I6[22], I7[22]);
	mux8to1 g23(Result[23], S, I0[23], I1[23], I2[23], I3[23], I4[23], I5[23], I6[23], I7[23]);
	mux8to1 g24(Result[24], S, I0[24], I1[24], I2[24], I3[24], I4[24], I5[24], I6[24], I7[24]);
	mux8to1 g25(Result[25], S, I0[25], I1[25], I2[25], I3[25], I4[25], I5[25], I6[25], I7[25]);
	mux8to1 g26(Result[26], S, I0[26], I1[26], I2[26], I3[26], I4[26], I5[26], I6[26], I7[26]);
	mux8to1 g27(Result[27], S, I0[27], I1[27], I2[27], I3[27], I4[27], I5[27], I6[27], I7[27]);
	mux8to1 g28(Result[28], S, I0[28], I1[28], I2[28], I3[28], I4[28], I5[28], I6[28], I7[28]);
	mux8to1 g29(Result[29], S, I0[29], I1[29], I2[29], I3[29], I4[29], I5[29], I6[29], I7[29]);
	mux8to1 g30(Result[30], S, I0[30], I1[30], I2[30], I3[30], I4[30], I5[30], I6[30], I7[30]);
	mux8to1 g31(Result[31], S, I0[31], I1[31], I2[31], I3[31], I4[31], I5[31], I6[31], I7[31]);


endmodule 