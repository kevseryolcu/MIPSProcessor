library verilog;
use verilog.vl_types.all;
entity genProp16bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end genProp16bit;
