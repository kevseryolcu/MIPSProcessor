library verilog;
use verilog.vl_types.all;
entity Adder32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end Adder32Bit;
