library verilog;
use verilog.vl_types.all;
entity and32Bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end and32Bit;
